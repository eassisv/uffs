library IEEE;

use IEEE.STD_LOGIC_1164.ALL;


entity mux4 is
    
Port ( SEL : in  STD_LOGIC;
           
       A   : in  STD_LOGIC;
        
       B   : in  STD_LOGIC;
         
       X   : out STD_LOGIC );

end mux4;



architecture comportamento of mux4 is
begin
    X <= A when (SEL = '1') else B;
end comportamento;


